import noc_params::*;

module circular_buffer #(
  parameter BUFFER_SIZE = VC_DEPTH;
)(
    input flit_t data_i,
    input read_i,
    input write_i,
    input rst,
    input clk,
    output flit_t data_o,
    output logic is_full,
    output logic is_empty
);

    localparam int POINTER_SIZE = $clog2(BUFFER_SIZE);

    flit_t memory[BUFFER_SIZE-1:0];

    logic [POINTER_SIZE-1:0] read_ptr;
    logic [POINTER_SIZE-1:0] write_ptr;

    logic [POINTER_SIZE-1:0] read_ptr_next;
    logic [POINTER_SIZE-1:0] write_ptr_next;

    logic [POINTER_SIZE:0] num_flits;
    logic [POINTER_SIZE:0] num_flits_next;

  	assign is_empty = (num_flits == 0);
  	assign is_full = (num_flits == BUFFER_SIZE);
    
    /*
    Sequential logic:
    - reset on the rising edge of the rst input;
    - when the write_i input is asserted on the rising edge of the clock,
      new data is added to the buffer
      or a simultaneous read is performed (i.e., the read_i input is asserted). Same for read_i.
    */
    always_ff@(posedge clk or posedge rst)
    begin
        if (rst)
        begin
            read_ptr    <= 0;
            write_ptr   <= 0;
            num_flits   <= 0;
          	data_o      <= 0;

        end
        else
        begin
            read_ptr    <= read_ptr_next;
            write_ptr   <= write_ptr_next;
            num_flits   <= num_flits_next;

          if (write_i)
                memory[write_ptr] <= data_i;
          
          if (read_i)
            	data_o <= memory[read_ptr];
        end
    end

    /*
    Combinational logic:
     FIFO contract:
	- read_i must only be asserted when is_empty == 0
	- write_i must only be asserted when is_full == 0
	- simultaneous read_i and write_i is allowed
	- FIFO does not perform internal legality checks
        * full and empty flags are eventually updated
        * read and write pointers are eventually incremented
        * the number of stored flits is updated
    - otherwise, the buffer next status doesn't change//
    */
    always_comb
    begin      
        unique if(read_i & ~write_i)
        begin: read_not_empty
            read_ptr_next = increase_ptr(read_ptr);
            write_ptr_next = write_ptr;
            num_flits_next = num_flits - 1;
        end
        else if(~read_i & write_i)
        begin: write_not_full
            read_ptr_next = read_ptr;
            write_ptr_next = increase_ptr(write_ptr);
            num_flits_next = num_flits + 1;
        end
        else if(read_i & write_i)
        begin: read_write_not_empty
            read_ptr_next = increase_ptr(read_ptr);
            write_ptr_next = increase_ptr(write_ptr);
            num_flits_next = num_flits;
        end
        else
        begin: do_nothing
            read_ptr_next = read_ptr;
            write_ptr_next = write_ptr;
            num_flits_next = num_flits;
        end
    end

    function logic [POINTER_SIZE-1:0] increase_ptr (input logic [POINTER_SIZE-1:0] ptr);
        if(ptr == BUFFER_SIZE-1)
            increase_ptr = 0;
        else
            increase_ptr = ptr+1;
    endfunction

endmodule
